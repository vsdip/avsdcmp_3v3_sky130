* SPICE3 file created from comparator.ext - technology: sky130A

.option scale=10000u

X0 VOUT a_305_n627# VDD w_n243_100# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=50
X1 VDD a_83_n114# a_198_n100# w_n243_100# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=600 l=50
X2 a_495_n214# a_198_n100# a_305_n627# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=5.20909e+06 ps=0 w=200 l=50
X3 a_83_n114# INP a_n86_n114# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=9 pd=98 as=1.06853e+09 ps=0 w=100 l=50
X4 VDD a_n208_n114# a_n208_n114# w_n243_100# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=8 ps=78 w=100 l=100
X5 GND VDD a_198_n100# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=1 as=0 ps=0 w=50 l=50
X6 a_181_n429# Ihyst GND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=1 as=0 ps=0 w=50 l=50
X7 GND EN a_495_n214# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=50
X8 VOUT a_305_n627# GND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=50
X9 a_n86_n114# INN a_n208_n114# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=100 l=50
X10 a_83_n114# a_198_n100# a_181_n429# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=50
X11 a_305_n627# a_198_n100# VDD w_n243_100# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=50
X12 a_83_n114# a_n208_n114# VDD w_n243_100# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=100 l=100
X13 a_181_n429# a_305_n627# a_n208_n114# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=200 l=50
X14 VDD EN a_305_n627# w_n243_100# sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=50
X15 Ihyst Ihyst GND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=8 pd=78 as=0 ps=0 w=50 l=50
X16 GND VDD a_n57_n429# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=9 ps=0 w=50 l=100
C0 GND a_305_n627# 2.06fF
C1 VDD SUB 6.17fF
C2 a_n208_n114# SUB 2.19fF
C3 a_198_n100# SUB 2.60fF
C4 w_n243_100# SUB 8.87fF
