**.subckt test_comparator
Ihyst VCC net4 0.8u
V1 VCC GND 3.3
V2 INN GND 1.235
V3 INP GND pwl 0 0.8 10u 1.8 20u 0.8 30u 1.8 40u 0.8 50u 1.8 60u 0.8 70u 1.8 80u 0.8 90u 1.8 100u
+ 0.8
XM3 net1 INN net2 GND sky130_fd_pr__nfet_03v3_nvt L=0.8 W=0.42
XM4 VDIFF INP net2 GND sky130_fd_pr__nfet_03v3_nvt L=0.8 W=0.42
XM8 net1 VOUT2 net3 GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 
XM9 VDIFF VOUT1 net3 GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 
XM5 net2 VCC GND GND sky130_fd_pr__nfet_03v3_nvt L=0.8 W=0.42 
XM2 VDIFF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 
XM1 net1 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 
XM12 VOUT2 VOUT1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 
XM10 VOUT1 VDIFF VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=6 
XM13 VOUT2 VOUT1 net5 GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=4  
XM11 VOUT1 VCC GND GND sky130_fd_pr__nfet_03v3_nvt L=0.8 W=0.42  
XM7 net3 net4 GND GND sky130_fd_pr__nfet_03v3_nvt L=0.8 W=0.42 
XM6 net4 net4 GND GND sky130_fd_pr__nfet_03v3_nvt L=0.6 W=0.42 
V4 EN GND 3.3
LOAD VOUT GND 10M m=1
XM14 VDIFF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 
XM15 net1 net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 
XM16 VOUT VOUT2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 
XM18 VOUT VOUT2 GND GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.42 
XM19 net5 EN GND GND sky130_fd_pr__nfet_03v3_nvt L=0.5 W=0.42 
XM22 VOUT2 EN VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 
**** begin user architecture code


.include ../Libs/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ../Libs/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
* Mismatch parameters
.include ../Libs/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ../Libs/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
*
* All models
.include ../Libs/models/all_mod.spice
*




.options savecurrents
.control
tran 10n 20u
# plot PLUS MINUS VDIFF V2nd VOUT
# plot net1 net2 net3
plot INP EN INN VOUT
plot VOUT vs INP-INN
.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
